SPICE3 Voltage meter

* Node 0 = GND
r1 1 2 1M
r2 2 0 100k
vdc 1 0 DC 12

.control
  * dispose of any 'save' statements from previous runs
  delete all
  dc vdc 0.5 24.0 0.5
  * draw a graph of the voltage vs time.
  plot  v(1),v(2)
  * print the voltage vs time
  print v(1),v(2)
.endc

.end
